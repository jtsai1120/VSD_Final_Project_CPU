
module Controller ();




endmodule